magic
tech gf180mcuD
timestamp 1755245820
<< nwell >>
rect -17 32 88 96
rect 25 31 75 32
<< nmos >>
rect -1 -7 5 10
rect 16 -7 22 10
rect 33 -7 39 10
rect 50 -7 56 10
rect 67 -7 73 10
<< pmos >>
rect 5 41 11 75
rect 16 41 22 75
rect 33 41 39 75
rect 50 41 56 75
rect 61 41 67 75
<< ndiff >>
rect -11 8 -1 10
rect -11 -5 -9 8
rect -4 -5 -1 8
rect -11 -7 -1 -5
rect 5 8 16 10
rect 5 0 8 8
rect 13 0 16 8
rect 5 -7 16 0
rect 22 8 33 10
rect 22 -5 25 8
rect 30 -5 33 8
rect 22 -7 33 -5
rect 39 8 50 10
rect 39 -5 42 8
rect 47 -5 50 8
rect 39 -7 50 -5
rect 56 3 67 10
rect 56 -5 59 3
rect 64 -5 67 3
rect 56 -7 67 -5
rect 73 8 83 10
rect 73 -5 76 8
rect 81 -5 83 8
rect 73 -7 83 -5
<< pdiff >>
rect -5 73 5 75
rect -5 43 -3 73
rect 2 43 5 73
rect -5 41 5 43
rect 11 41 16 75
rect 22 73 33 75
rect 22 43 25 73
rect 30 43 33 73
rect 22 41 33 43
rect 39 73 50 75
rect 39 43 42 73
rect 47 43 50 73
rect 39 41 50 43
rect 56 41 61 75
rect 67 73 77 75
rect 67 43 70 73
rect 75 43 77 73
rect 67 41 77 43
<< ndiffc >>
rect -9 -5 -4 8
rect 8 0 13 8
rect 25 -5 30 8
rect 42 -5 47 8
rect 59 -5 64 3
rect 76 -5 81 8
<< pdiffc >>
rect -3 43 2 73
rect 25 43 30 73
rect 42 43 47 73
rect 70 43 75 73
<< psubdiff >>
rect -14 -19 1 -17
rect -14 -24 -9 -19
rect -4 -24 1 -19
rect -14 -26 1 -24
rect 7 -19 22 -17
rect 7 -24 12 -19
rect 17 -24 22 -19
rect 7 -26 22 -24
rect 28 -19 43 -17
rect 28 -24 33 -19
rect 38 -24 43 -19
rect 28 -26 43 -24
rect 49 -19 64 -17
rect 49 -24 54 -19
rect 59 -24 64 -19
rect 49 -26 64 -24
rect 70 -19 85 -17
rect 70 -24 75 -19
rect 80 -24 85 -19
rect 70 -26 85 -24
<< nsubdiff >>
rect -14 89 1 91
rect -14 84 -9 89
rect -4 84 1 89
rect -14 82 1 84
rect 7 89 22 91
rect 7 84 12 89
rect 17 84 22 89
rect 7 82 22 84
rect 28 89 43 91
rect 28 84 33 89
rect 38 84 43 89
rect 28 82 43 84
rect 49 89 64 91
rect 49 84 54 89
rect 59 84 64 89
rect 49 82 64 84
rect 70 89 85 91
rect 70 84 75 89
rect 80 84 85 89
rect 70 82 85 84
<< psubdiffcont >>
rect -9 -24 -4 -19
rect 12 -24 17 -19
rect 33 -24 38 -19
rect 54 -24 59 -19
rect 75 -24 80 -19
<< nsubdiffcont >>
rect -9 84 -4 89
rect 12 84 17 89
rect 33 84 38 89
rect 54 84 59 89
rect 75 84 80 89
<< polysilicon >>
rect 5 75 11 80
rect 16 75 22 80
rect 33 75 39 80
rect 50 75 56 80
rect 61 75 67 80
rect 5 39 11 41
rect -1 33 11 39
rect -1 25 5 33
rect 16 25 22 41
rect 33 28 39 41
rect 50 28 56 41
rect 61 39 67 41
rect 61 33 73 39
rect 67 28 73 33
rect 34 26 44 28
rect -7 23 3 25
rect -7 17 -5 23
rect 1 17 3 23
rect -7 15 3 17
rect 18 23 28 25
rect 18 17 20 23
rect 26 17 28 23
rect 34 20 36 26
rect 42 20 44 26
rect 34 18 44 20
rect 50 26 60 28
rect 50 20 52 26
rect 58 20 60 26
rect 50 18 60 20
rect 66 26 76 28
rect 66 20 68 26
rect 74 20 76 26
rect 66 18 76 20
rect 18 15 28 17
rect -1 10 5 15
rect 16 10 22 15
rect 33 10 39 18
rect 50 10 56 18
rect 67 10 73 18
rect -1 -12 5 -7
rect 16 -12 22 -7
rect 33 -12 39 -7
rect 50 -12 56 -7
rect 67 -12 73 -7
<< polycontact >>
rect -5 17 1 23
rect 20 17 26 23
rect 36 20 42 26
rect 52 20 58 26
rect 68 20 74 26
<< metal1 >>
rect -17 89 88 96
rect -17 84 -9 89
rect -4 84 12 89
rect 17 84 33 89
rect 38 84 54 89
rect 59 84 75 89
rect 80 84 88 89
rect -17 82 88 84
rect -3 73 2 82
rect -3 41 2 43
rect 25 73 30 75
rect 25 36 30 43
rect 42 73 47 82
rect 42 41 47 43
rect 70 73 75 75
rect 70 40 75 43
rect 70 36 77 40
rect 8 34 77 36
rect 83 34 85 40
rect 8 31 75 34
rect -7 17 -5 23
rect 1 17 3 23
rect -9 8 -4 10
rect 8 8 13 31
rect 18 17 20 23
rect 26 17 28 23
rect 34 20 36 26
rect 42 20 44 26
rect 50 20 52 26
rect 58 20 60 26
rect 66 20 68 26
rect 74 20 76 26
rect 42 10 81 15
rect 8 -2 13 0
rect 25 8 30 10
rect -9 -7 -4 -5
rect 25 -7 30 -5
rect 42 8 47 10
rect 76 8 81 10
rect 42 -7 47 -5
rect 59 3 64 5
rect -9 -12 30 -7
rect 59 -17 64 -5
rect 76 -7 81 -5
rect -17 -19 88 -17
rect -17 -24 -9 -19
rect -4 -24 12 -19
rect 17 -24 33 -19
rect 38 -24 54 -19
rect 59 -24 75 -19
rect 80 -24 88 -19
rect -17 -31 88 -24
<< via1 >>
rect 77 34 83 40
rect -5 17 1 23
rect 20 17 26 23
rect 36 20 42 26
rect 52 20 58 26
rect 68 20 74 26
<< metal2 >>
rect 76 40 84 41
rect 76 34 77 40
rect 83 34 84 40
rect 76 33 84 34
rect 34 26 44 27
rect -7 23 3 24
rect -7 17 -5 23
rect 1 17 3 23
rect -7 16 3 17
rect 18 23 28 24
rect 18 17 20 23
rect 26 17 28 23
rect 34 20 36 26
rect 42 20 44 26
rect 34 19 44 20
rect 50 26 60 27
rect 50 20 52 26
rect 58 20 60 26
rect 50 19 60 20
rect 66 26 76 27
rect 66 20 68 26
rect 74 20 76 26
rect 66 19 76 20
rect 18 16 28 17
<< labels >>
rlabel metal2 -5 17 1 23 1 A0
rlabel metal2 20 17 26 23 1 A1
rlabel metal2 36 20 42 26 1 C
rlabel metal2 52 20 58 26 1 B0
rlabel metal2 68 20 74 26 1 B1
rlabel via1 77 34 83 40 1 Y
rlabel nsubdiffcont -9 84 -4 89 1 vdd
rlabel psubdiffcont -9 -24 -4 -19 1 vss
<< end >>
