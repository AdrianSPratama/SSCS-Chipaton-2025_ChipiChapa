* NGSPICE file created from gf180mcu_gp9t3v3__aoi221_1.ext - technology: gf180mcuD

**.subckt gf180mcu_gp9t3v3__aoi221_1 A0 A1 B0 B1 C Y vdd vss
X0 a_30_670# B0 vdd vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1 Y A1 a_530_670# vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X2 a_250_160# B1 vss vss nfet_03v3 ad=0.10625p pd=1.1u as=0.425p ps=2.7u w=0.85u l=0.3u
X3 vss C Y vss nfet_03v3 ad=0.27625p pd=1.5u as=0.27625p ps=1.5u w=0.85u l=0.3u
X4 a_530_670# A0 Y vdd pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 Y A0 a_740_160# vss nfet_03v3 ad=0.425p pd=2.7u as=0.10625p ps=1.1u w=0.85u l=0.3u
X6 vdd B1 a_30_670# vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X7 Y B0 a_250_160# vss nfet_03v3 ad=0.27625p pd=1.5u as=0.10625p ps=1.1u w=0.85u l=0.3u
X8 a_740_160# A1 vss vss nfet_03v3 ad=0.10625p pd=1.1u as=0.27625p ps=1.5u w=0.85u l=0.3u
X9 a_530_670# C a_30_670# vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
**.ends

