VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_gp9t3v3_oai211_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_gp9t3v3_oai211_1 ;
  ORIGIN 3.000 2.850 ;
  SIZE 4.450 BY 6.350 ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT -2.600 0.000 -2.100 0.300 ;
      LAYER Metal2 ;
        RECT -2.600 -0.050 -2.100 0.350 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT -1.500 0.000 -1.000 0.300 ;
      LAYER Metal2 ;
        RECT -1.500 -0.050 -1.000 0.350 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT -0.700 0.000 -0.200 0.300 ;
      LAYER Metal2 ;
        RECT -0.700 -0.050 -0.200 0.350 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.100 0.000 0.600 0.300 ;
      LAYER Metal2 ;
        RECT 0.100 -0.050 0.600 0.350 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.210000 ;
    PORT
      LAYER Metal1 ;
        RECT -1.050 1.100 -0.800 1.850 ;
        RECT 0.650 1.100 0.900 1.850 ;
        RECT -1.050 0.850 0.900 1.100 ;
        RECT 0.650 0.800 0.900 0.850 ;
        RECT 0.650 0.550 1.200 0.800 ;
        RECT 0.950 -0.300 1.200 0.550 ;
        RECT 0.800 -0.650 1.200 -0.300 ;
        RECT 0.650 -0.950 1.200 -0.650 ;
        RECT 0.650 -1.650 0.900 -0.950 ;
      LAYER Metal2 ;
        RECT 0.800 -0.700 1.200 -0.300 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -3.000 0.300 1.450 3.500 ;
      LAYER Metal1 ;
        RECT -3.000 2.800 1.450 3.500 ;
        RECT -2.450 1.500 -2.200 2.800 ;
        RECT -0.200 1.500 0.050 2.800 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT -1.600 -2.150 -1.350 -1.200 ;
        RECT -3.000 -2.850 1.450 -2.150 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT -2.450 -0.950 -0.500 -0.700 ;
        RECT -2.450 -1.650 -2.200 -0.950 ;
        RECT -0.750 -1.650 -0.500 -0.950 ;
  END
END gf180mcu_gp9t3v3_oai211_1
END LIBRARY

