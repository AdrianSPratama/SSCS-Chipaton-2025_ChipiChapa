VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_gp9t3v3_oai221_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_gp9t3v3_oai221_1 ;
  ORIGIN 0.850 1.550 ;
  SIZE 5.250 BY 6.350 ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT -0.350 0.850 0.150 1.150 ;
      LAYER Metal2 ;
        RECT -0.350 0.800 0.150 1.200 ;
    END
  END A0
  PIN A1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 0.850 1.400 1.150 ;
      LAYER Metal2 ;
        RECT 0.900 0.800 1.400 1.200 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.500 1.000 3.000 1.300 ;
      LAYER Metal2 ;
        RECT 2.500 0.950 3.000 1.350 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.300 1.000 3.800 1.300 ;
      LAYER Metal2 ;
        RECT 3.300 0.950 3.800 1.350 ;
    END
  END B1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.700 1.000 2.200 1.300 ;
      LAYER Metal2 ;
        RECT 1.700 0.950 2.200 1.350 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.252500 ;
    PORT
      LAYER Metal1 ;
        RECT 1.250 1.800 1.500 3.750 ;
        RECT 3.500 2.000 3.750 3.750 ;
        RECT 3.500 1.800 4.250 2.000 ;
        RECT 0.400 1.700 4.250 1.800 ;
        RECT 0.400 1.550 3.750 1.700 ;
        RECT 0.400 -0.100 0.650 1.550 ;
      LAYER Metal2 ;
        RECT 3.800 1.650 4.200 2.050 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -0.850 1.600 4.400 4.800 ;
        RECT 1.250 1.550 3.750 1.600 ;
      LAYER Metal1 ;
        RECT -0.850 4.100 4.400 4.800 ;
        RECT -0.150 2.050 0.100 4.100 ;
        RECT 2.100 2.050 2.350 4.100 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.950 -0.850 3.200 0.250 ;
        RECT -0.850 -1.550 4.400 -0.850 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 2.100 0.500 4.050 0.750 ;
        RECT -0.450 -0.350 -0.200 0.500 ;
        RECT 1.250 -0.350 1.500 0.500 ;
        RECT 2.100 -0.350 2.350 0.500 ;
        RECT 3.800 -0.350 4.050 0.500 ;
        RECT -0.450 -0.600 1.500 -0.350 ;
  END
END gf180mcu_gp9t3v3_oai221_1
END LIBRARY

