* SPICE3 file created from gf180mcu_gp9t3v3__aoi221_1.2.ext - technology: gf180mcuD

.option scale=5n

X0 a_30_670# B0.t0 vdd.t1 vdd.t0 pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
X1 Y.t1 A1.t0 a_530_670# vdd.t2 pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
X2 a_250_160# B1.t0 vss.t7 vss.t6 nfet_03v3 ad=4.25n pd=0.22m as=17n ps=0.54m w=170 l=60
X3 vss.t5 C.t0 Y.t3 vss.t4 nfet_03v3 ad=11.05n pd=0.3m as=11.05n ps=0.3m w=170 l=60
X4 a_530_670# A0.t0 Y.t4 vdd.t6 pfet_03v3 ad=34n pd=0.88m as=18.7n ps=0.45m w=340 l=60
X5 Y.t2 A0.t1 a_740_160# vss.t3 nfet_03v3 ad=17n pd=0.54m as=4.25n ps=0.22m w=170 l=60
X6 vdd.t5 B1.t1 a_30_670# vdd.t4 pfet_03v3 ad=18.7n pd=0.45m as=34n ps=0.88m w=340 l=60
X7 Y.t0 B0.t1 a_250_160# vss.t0 nfet_03v3 ad=11.05n pd=0.3m as=4.25n ps=0.22m w=170 l=60
X8 a_740_160# A1.t1 vss.t2 vss.t1 nfet_03v3 ad=4.25n pd=0.22m as=11.05n ps=0.3m w=170 l=60
X9 a_530_670# C.t1 a_30_670# vdd.t3 pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
C0 Y a_530_670# 0.10318f
C1 A1 a_530_670# 0.03341f
C2 Y A1 0.21331f
C3 B0 vdd 0.10252f
C4 a_740_160# Y 0.0043f
C5 B0 a_530_670# 0.00134f
C6 Y B0 0.00974f
C7 B0 A1 0
C8 vdd A0 0.12702f
C9 C vdd 0.10597f
C10 A0 a_530_670# 0.04623f
C11 vdd B1 0.10787f
C12 vdd a_30_670# 0.17787f
C13 C a_530_670# 0.00502f
C14 a_30_670# a_530_670# 0.02429f
C15 Y A0 0.21193f
C16 A0 A1 0.07085f
C17 Y C 0.13459f
C18 C A1 0.11332f
C19 Y B1 0.00897f
C20 Y a_30_670# 0.04804f
C21 A1 B1 0
C22 A1 a_30_670# 0.00307f
C23 a_250_160# Y 0
C24 B0 A0 0
C25 C B0 0.10697f
C26 B0 B1 0.11641f
C27 B0 a_30_670# 0.1005f
C28 a_250_160# B0 0.00221f
C29 C A0 0
C30 vdd a_530_670# 0.26686f
C31 A0 B1 0
C32 A0 a_30_670# 0
C33 C B1 0
C34 C a_30_670# 0.01213f
C35 Y vdd 0.02607f
C36 B1 a_30_670# 0.08494f
C37 vdd A1 0.08965f
C38 a_250_160# a_30_670# 0
R0 B0 B0.t0 50.4922
R1 B0.t1 B0.n0 39.5422
R2 B0 B0.t1 20.0755
R3 vdd.t3 vdd.t2 265.625
R4 vdd.n3 vdd.t0 257.812
R5 vdd.t4 vdd.n6 195.312
R6 vdd.n7 vdd.t4 145.413
R7 vdd.n2 vdd.t6 77.536
R8 vdd.n6 vdd.t0 70.313
R9 vdd.t2 vdd.n2 62.2079
R10 vdd.n4 vdd.n3 12.6005
R11 vdd.n6 vdd.n5 12.6005
R12 vdd.n3 vdd.t3 7.813
R13 vdd.n4 vdd.n2 4.76743
R14 vdd.n1 vdd.n0 2.88873
R15 vdd.n0 vdd.t1 1.13285
R16 vdd.n0 vdd.t5 1.13285
R17 vdd.n5 vdd.n4 0.1355
R18 vdd.n7 vdd.n1 0.109786
R19 vdd vdd.n7 0.0872857
R20 vdd.n5 vdd.n1 0.0262143
R21 A1 A1.t0 47.4505
R22 A1 A1.t1 23.7255
R23 Y.n3 Y.t2 8.59974
R24 Y.n2 Y.n1 7.2005
R25 Y Y.n4 4.54005
R26 Y.n2 Y.n0 3.15473
R27 Y.n1 Y.t3 2.77991
R28 Y.n1 Y.t0 2.03874
R29 Y.n0 Y.t4 1.13285
R30 Y.n0 Y.t1 1.13285
R31 Y.n3 Y.n2 0.1535
R32 Y.n4 Y.n3 0.1115
R33 B1 B1.t1 40.1505
R34 B1.n1 B1.t0 19.4672
R35 B1.n1 B1.n0 8.92272
R36 B1 B1.n1 8.51717
R37 vss.t4 vss.n4 954.365
R38 vss.n5 vss.t0 851.191
R39 vss.n9 vss.t6 758.417
R40 vss.t3 vss.t1 567.461
R41 vss.n3 vss.t3 500.615
R42 vss.t6 vss.n8 335.317
R43 vss.n8 vss.t0 232.143
R44 vss.n5 vss.t4 128.969
R45 vss.n4 vss.t1 25.7941
R46 vss.n4 vss.n3 10.4005
R47 vss.n6 vss.n5 10.4005
R48 vss.n8 vss.n7 10.4005
R49 vss.n0 vss.t7 8.60874
R50 vss.n2 vss.n1 6.5615
R51 vss.n1 vss.t5 2.77991
R52 vss.n1 vss.t2 2.03874
R53 vss.n7 vss.n6 0.1355
R54 vss.n7 vss.n0 0.0969286
R55 vss vss.n9 0.0872857
R56 vss.n6 vss.n2 0.0840714
R57 vss.n3 vss.n2 0.0519286
R58 vss.n9 vss.n0 0.0390714
R59 C C.t1 47.4505
R60 C C.t0 23.7255
R61 A0 A0.t0 52.9498
R62 A0.t1 A0.n0 41.9755
R63 A0 A0.t1 22.5088
C39 Y vss 0.57547f
C40 A0 vss 0.37725f
C41 A1 vss 0.29923f
C42 C vss 0.29661f
C43 B0 vss 0.30231f
C44 B1 vss 0.43242f
C45 vdd vss 2.41757f
C46 a_740_160# vss 0.00366f
C47 a_250_160# vss 0.00366f 
C48 a_530_670# vss 0.05393f 
C49 a_30_670# vss 0.09822f
