* SPICE3 file created from gf180mcu_gp9t3v3_oai211_1.ext - technology: gf180mcuD
.subckt gf180mcu_gp9t3v3_oai211_1 vdd Y A0 A1 B C vss
X0 Y C vdd vdd pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1 a_n350_150# A0 vdd vdd pfet_03v3 ad=0.2125p pd=1.95u as=0.85p ps=4.4u w=1.7u l=0.3u
X2 a_n510_n360# A1 vss vss nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3 Y C a_n10_n360# vss nfet_03v3 ad=0.425p pd=2.7u as=0.10625p ps=1.1u w=0.85u l=0.3u
X4 Y A1 a_n350_150# vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.2125p ps=1.95u w=1.7u l=0.3u
X5 vdd B Y vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X6 vss A0 a_n510_n360# vss nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X7 a_n10_n360# B a_n510_n360# vss nfet_03v3 ad=0.10625p pd=1.1u as=0.23375p ps=1.4u w=0.85u l=0.3u
C0 C Y 0.1582f
C1 a_n510_n360# vdd 0.01219f
C2 A0 vdd 0.11214f
C3 A1 vdd 0.1015f
C4 a_n510_n360# C 0.00287f
C5 a_n10_n360# C 0
C6 vdd B 0.10701f
C7 Y a_n350_150# 0.00202f
C8 C B 0.16806f
C9 a_n510_n360# a_n350_150# 0.00253f
C10 a_n510_n360# Y 0.04443f
C11 a_n10_n360# Y 0.00215f
C12 C vdd 0.10654f
C13 A0 Y 0.00421f
C14 A1 Y 0.01623f
C15 a_n10_n360# a_n510_n360# 0.00112f
C16 A0 a_n510_n360# 0.07815f
C17 A1 a_n510_n360# 0.07761f
C18 A1 A0 0.17698f
C19 Y B 0.06331f
C20 a_n510_n360# B 0.02683f
C21 vdd a_n350_150# 0.00727f
C22 A1 B 0.14798f
C23 Y vdd 0.24175f
C24 Y vss 0.31362f
C25 C vss 0.3293f
C26 B vss 0.28763f
C27 A1 vss 0.28567f
C28 A0 vss 0.34649f
C29 vdd vss 1.96279f
C30 a_n10_n360# vss 0.00315f
C31 a_n510_n360# vss 0.30297f
.ends