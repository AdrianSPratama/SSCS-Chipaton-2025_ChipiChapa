VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_gp9t3v3__aoi221_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_gp9t3v3__aoi221_1 ;
  ORIGIN 0.300 0.250 ;
  SIZE 5.600 BY 6.350 ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.350 2.700 4.850 3.000 ;
      LAYER Metal2 ;
        RECT 4.350 2.650 4.850 3.050 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 2.300 3.600 2.600 ;
      LAYER Metal2 ;
        RECT 3.100 2.250 3.600 2.650 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.300 2.250 1.800 2.550 ;
      LAYER Metal2 ;
        RECT 1.300 2.200 1.800 2.600 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.450 2.100 0.950 2.400 ;
      LAYER Metal2 ;
        RECT 0.450 2.050 0.950 2.450 ;
    END
  END B1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.200 2.300 2.700 2.600 ;
      LAYER Metal2 ;
        RECT 2.200 2.250 2.700 2.650 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.912500 ;
    PORT
      LAYER Metal1 ;
        RECT 3.650 3.100 3.900 4.300 ;
        RECT 3.650 2.850 4.100 3.100 ;
        RECT 3.850 2.050 4.100 2.850 ;
        RECT 4.400 2.050 5.050 2.300 ;
        RECT 1.950 2.000 5.050 2.050 ;
        RECT 1.950 1.800 4.650 2.000 ;
        RECT 1.950 0.800 2.200 1.800 ;
        RECT 4.400 0.800 4.650 1.800 ;
      LAYER Metal2 ;
        RECT 4.500 1.950 5.050 2.350 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -0.300 2.900 5.300 6.100 ;
      LAYER Metal1 ;
        RECT -0.300 5.400 5.300 6.100 ;
        RECT 1.100 3.950 1.350 5.400 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.450 0.800 1.600 ;
        RECT 3.000 0.450 3.250 1.550 ;
        RECT -0.300 -0.250 5.300 0.450 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 2.800 4.750 4.750 5.000 ;
        RECT 0.250 3.150 0.500 4.300 ;
        RECT 1.950 3.150 2.200 4.300 ;
        RECT 2.800 4.050 3.050 4.750 ;
        RECT 4.500 4.050 4.750 4.750 ;
        RECT 0.250 2.900 2.200 3.150 ;
  END
END gf180mcu_gp9t3v3__aoi221_1
END LIBRARY

