* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3_aoi211_1.ext - technology: gf180mcuD

.option scale=5n

X0 a_70_30# A1 vss vss nfet_03v3 ad=9.35n pd=0.28m as=17n ps=0.54m w=170 l=60
X1 vdd A1 a_n90_540# vdd pfet_03v3 ad=18.7n pd=0.45m as=34n ps=0.88m w=340 l=60
X2 Y C a_410_540# vdd pfet_03v3 ad=34n pd=0.88m as=8.5n ps=0.39m w=340 l=60
X3 Y C vss vss nfet_03v3 ad=17n pd=0.54m as=9.35n ps=0.28m w=170 l=60
X4 a_n90_540# A0 vdd vdd pfet_03v3 ad=18.7n pd=0.45m as=18.7n ps=0.45m w=340 l=60
X5 vss B Y vss nfet_03v3 ad=9.35n pd=0.28m as=9.35n ps=0.28m w=170 l=60
X6 Y A0 a_70_30# vss nfet_03v3 ad=9.35n pd=0.28m as=9.35n ps=0.28m w=170 l=60
X7 a_410_540# B a_n90_540# vdd pfet_03v3 ad=8.5n pd=0.39m as=18.7n ps=0.45m w=340 l=60
C0 vdd C 0.10468f
C1 Y a_70_30# 0.00155f
C2 B Y 0.107f
C3 B vdd 0.09771f
C4 Y A0 0.00888f
C5 C a_n90_540# 0.00365f
C6 A0 vdd 0.10437f
C7 Y A1 0.00361f
C8 vdd A1 0.1078f
C9 a_70_30# a_n90_540# 0.00184f
C10 B a_n90_540# 0.01634f
C11 B C 0.17532f
C12 A0 a_n90_540# 0.05759f
C13 a_n90_540# A1 0.0598f
C14 Y a_410_540# 0.00464f
C15 a_410_540# vdd 0.00522f
C16 A0 a_70_30# 0.00209f
C17 B A0 0.14253f
C18 Y vdd 0.07048f
C19 a_410_540# a_n90_540# 0.00262f
C20 A0 A1 0.1279f
C21 Y a_n90_540# 0.04331f
C22 vdd a_n90_540# 0.24256f
C23 Y C 0.22754f
C24 Y vss 0.54509f
C25 C vss 0.33792f
C26 B vss 0.28193f
C27 A0 vss 0.29139f
C28 A1 vss 0.36819f
C29 vdd vss 1.92733f
C30 a_70_30# vss 0.00844f **FLOATING
C31 a_n90_540# vss 0.09099f **FLOATING
