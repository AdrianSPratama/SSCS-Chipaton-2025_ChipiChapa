magic
tech gf180mcuD
timestamp 1754635369
<< nwell >>
rect -6 44 106 122
<< nmos >>
rect 19 15 25 35
rect 30 15 36 35
rect 49 20 55 30
rect 68 15 74 35
rect 79 15 85 35
<< pmos >>
rect 13 57 19 102
rect 30 57 36 102
rect 47 57 53 102
rect 64 57 70 102
rect 81 57 87 102
<< ndiff >>
rect 9 29 19 35
rect 9 17 11 29
rect 16 17 19 29
rect 9 15 19 17
rect 25 15 30 35
rect 36 33 47 35
rect 36 21 39 33
rect 44 30 47 33
rect 57 30 68 35
rect 44 21 49 30
rect 36 20 49 21
rect 55 29 68 30
rect 55 20 60 29
rect 36 15 47 20
rect 57 17 60 20
rect 65 17 68 29
rect 57 15 68 17
rect 74 15 79 35
rect 85 33 95 35
rect 85 21 88 33
rect 93 21 95 33
rect 85 15 95 21
<< pdiff >>
rect 3 75 13 102
rect 3 70 5 75
rect 10 70 13 75
rect 3 65 13 70
rect 3 60 5 65
rect 10 60 13 65
rect 3 57 13 60
rect 19 98 30 102
rect 19 93 22 98
rect 27 93 30 98
rect 19 88 30 93
rect 19 83 22 88
rect 27 83 30 88
rect 19 57 30 83
rect 36 75 47 102
rect 36 70 39 75
rect 44 70 47 75
rect 36 65 47 70
rect 36 60 39 65
rect 44 60 47 65
rect 36 57 47 60
rect 53 99 64 102
rect 53 94 56 99
rect 61 94 64 99
rect 53 89 64 94
rect 53 84 56 89
rect 61 84 64 89
rect 53 57 64 84
rect 70 75 81 102
rect 70 70 73 75
rect 78 70 81 75
rect 70 65 81 70
rect 70 60 73 65
rect 78 60 81 65
rect 70 57 81 60
rect 87 99 97 102
rect 87 94 90 99
rect 95 94 97 99
rect 87 89 97 94
rect 87 84 90 89
rect 95 84 97 89
rect 87 57 97 84
<< ndiffc >>
rect 11 17 16 29
rect 39 21 44 33
rect 60 17 65 29
rect 88 21 93 33
<< pdiffc >>
rect 5 70 10 75
rect 5 60 10 65
rect 22 93 27 98
rect 22 83 27 88
rect 39 70 44 75
rect 39 60 44 65
rect 56 94 61 99
rect 56 84 61 89
rect 73 70 78 75
rect 73 60 78 65
rect 90 94 95 99
rect 90 84 95 89
<< psubdiff >>
rect 0 5 15 7
rect 0 0 4 5
rect 9 0 15 5
rect 0 -2 15 0
rect 21 5 36 7
rect 21 0 26 5
rect 31 0 36 5
rect 21 -2 36 0
rect 42 5 57 7
rect 42 0 47 5
rect 52 0 57 5
rect 42 -2 57 0
rect 63 5 78 7
rect 63 0 68 5
rect 73 0 78 5
rect 63 -2 78 0
rect 84 5 99 7
rect 84 0 89 5
rect 94 0 99 5
rect 84 -2 99 0
<< nsubdiff >>
rect 3 117 18 119
rect 3 112 8 117
rect 13 112 18 117
rect 3 110 18 112
rect 24 117 39 119
rect 24 112 29 117
rect 34 112 39 117
rect 24 110 39 112
rect 45 117 60 119
rect 45 112 50 117
rect 55 112 60 117
rect 45 110 60 112
rect 66 117 81 119
rect 66 112 71 117
rect 76 112 81 117
rect 66 110 81 112
<< psubdiffcont >>
rect 4 0 9 5
rect 26 0 31 5
rect 47 0 52 5
rect 68 0 73 5
rect 89 0 94 5
<< nsubdiffcont >>
rect 8 112 13 117
rect 29 112 34 117
rect 50 112 55 117
rect 71 112 76 117
<< polysilicon >>
rect 13 102 19 107
rect 30 102 36 107
rect 47 102 53 107
rect 64 102 70 107
rect 81 102 87 107
rect 13 52 19 57
rect 30 55 36 57
rect 25 53 36 55
rect 47 54 53 57
rect 64 54 70 57
rect 81 55 87 57
rect 13 50 17 52
rect 8 47 17 50
rect 8 42 10 47
rect 15 42 17 47
rect 25 48 29 53
rect 34 48 36 53
rect 25 46 36 48
rect 8 41 17 42
rect 8 37 25 41
rect 32 40 36 46
rect 43 52 54 54
rect 43 47 47 52
rect 52 47 54 52
rect 61 52 72 54
rect 61 47 65 52
rect 70 47 72 52
rect 81 52 96 55
rect 81 51 89 52
rect 43 45 55 47
rect 61 45 72 47
rect 86 47 89 51
rect 94 47 96 52
rect 86 45 96 47
rect 19 35 25 37
rect 30 35 36 40
rect 51 35 55 45
rect 68 40 72 45
rect 81 41 96 45
rect 81 40 85 41
rect 68 35 74 40
rect 79 35 85 40
rect 49 30 55 35
rect 49 15 55 20
rect 19 10 25 15
rect 30 10 36 15
rect 68 10 74 15
rect 79 10 85 15
<< polycontact >>
rect 10 42 15 47
rect 29 48 34 53
rect 47 47 52 52
rect 65 47 70 52
rect 89 47 94 52
<< metal1 >>
rect -6 117 106 122
rect -6 112 8 117
rect 13 112 29 117
rect 34 112 50 117
rect 55 112 71 117
rect 76 112 106 117
rect -6 108 106 112
rect 22 98 27 108
rect 22 88 27 93
rect 22 80 27 83
rect 56 99 95 101
rect 61 96 90 99
rect 56 89 61 94
rect 56 82 61 84
rect 90 89 95 94
rect 90 82 95 84
rect 5 75 10 77
rect 5 65 10 70
rect 39 75 44 77
rect 39 65 44 70
rect 10 60 39 63
rect 5 58 44 60
rect 73 75 78 77
rect 73 65 78 70
rect 78 60 82 62
rect 73 57 82 60
rect 8 48 17 49
rect 4 42 9 48
rect 15 42 17 48
rect 23 47 28 53
rect 34 47 36 53
rect 41 46 46 52
rect 52 46 54 52
rect 59 46 64 52
rect 70 46 72 52
rect 8 41 17 42
rect 77 41 82 57
rect 87 46 89 52
rect 95 46 100 52
rect 39 36 93 41
rect 39 33 44 36
rect 11 29 16 31
rect 88 33 93 36
rect 39 19 44 21
rect 60 29 65 31
rect 11 9 16 17
rect 88 19 93 21
rect 60 9 65 17
rect -6 5 106 9
rect -6 0 4 5
rect 9 0 26 5
rect 31 0 47 5
rect 52 0 68 5
rect 73 0 89 5
rect 94 0 106 5
rect -6 -5 106 0
<< via1 >>
rect 9 47 15 48
rect 9 42 10 47
rect 10 42 15 47
rect 28 48 29 53
rect 29 48 34 53
rect 28 47 34 48
rect 46 47 47 52
rect 47 47 52 52
rect 46 46 52 47
rect 64 47 65 52
rect 65 47 70 52
rect 64 46 70 47
rect 89 47 94 52
rect 94 47 95 52
rect 89 46 95 47
<< metal2 >>
rect 25 53 36 54
rect 6 48 17 49
rect 6 42 9 48
rect 15 42 17 48
rect 25 47 28 53
rect 34 47 36 53
rect 25 46 36 47
rect 43 52 54 53
rect 43 46 46 52
rect 52 46 54 52
rect 43 45 54 46
rect 61 52 72 53
rect 61 46 64 52
rect 70 46 72 52
rect 61 45 72 46
rect 87 52 98 53
rect 87 46 89 52
rect 95 46 98 52
rect 87 45 98 46
rect 6 41 17 42
<< labels >>
rlabel metal1 -6 114 -6 114 3 vdd
rlabel metal1 -6 1 -6 1 3 vss
rlabel polysilicon 25 41 25 41 1 B1
rlabel polysilicon 36 40 36 40 1 B0
rlabel polysilicon 51 42 51 42 1 C
rlabel polysilicon 68 42 68 42 1 A1
rlabel polysilicon 96 41 96 41 1 A0
<< end >>
