magic
tech gf180mcuD
timestamp 1755145353
<< nwell >>
rect -60 6 29 70
<< nmos >>
rect -41 -36 -35 -19
rect -24 -36 -18 -19
rect -7 -36 -1 -19
rect 4 -36 10 -19
<< pmos >>
rect -41 15 -35 49
rect -30 15 -24 49
rect -13 15 -7 49
rect 4 15 10 49
<< ndiff >>
rect -51 -23 -41 -19
rect -51 -31 -49 -23
rect -44 -31 -41 -23
rect -51 -36 -41 -31
rect -35 -26 -24 -19
rect -35 -34 -32 -26
rect -27 -34 -24 -26
rect -35 -36 -24 -34
rect -18 -23 -7 -19
rect -18 -31 -15 -23
rect -10 -31 -7 -23
rect -18 -36 -7 -31
rect -1 -36 4 -19
rect 10 -23 20 -19
rect 10 -31 13 -23
rect 18 -31 20 -23
rect 10 -36 20 -31
<< pdiff >>
rect -51 47 -41 49
rect -51 42 -49 47
rect -44 42 -41 47
rect -51 37 -41 42
rect -51 32 -49 37
rect -44 32 -41 37
rect -51 15 -41 32
rect -35 15 -30 49
rect -24 34 -13 49
rect -24 29 -21 34
rect -16 29 -13 34
rect -24 24 -13 29
rect -24 19 -21 24
rect -16 19 -13 24
rect -24 15 -13 19
rect -7 47 4 49
rect -7 42 -4 47
rect 1 42 4 47
rect -7 37 4 42
rect -7 32 -4 37
rect 1 32 4 37
rect -7 15 4 32
rect 10 34 20 49
rect 10 29 13 34
rect 18 29 20 34
rect 10 24 20 29
rect 10 19 13 24
rect 18 19 20 24
rect 10 15 20 19
<< ndiffc >>
rect -49 -31 -44 -23
rect -32 -34 -27 -26
rect -15 -31 -10 -23
rect 13 -31 18 -23
<< pdiffc >>
rect -49 42 -44 47
rect -49 32 -44 37
rect -21 29 -16 34
rect -21 19 -16 24
rect -4 42 1 47
rect -4 32 1 37
rect 13 29 18 34
rect 13 19 18 24
<< psubdiff >>
rect -54 -45 -39 -43
rect -54 -50 -49 -45
rect -44 -50 -39 -45
rect -54 -52 -39 -50
rect -33 -45 -18 -43
rect -33 -50 -28 -45
rect -23 -50 -18 -45
rect -33 -52 -18 -50
rect -12 -45 3 -43
rect -12 -50 -7 -45
rect -2 -50 3 -45
rect -12 -52 3 -50
rect 9 -45 24 -43
rect 9 -50 14 -45
rect 19 -50 24 -45
rect 9 -52 24 -50
<< nsubdiff >>
rect -54 63 -39 65
rect -54 58 -49 63
rect -44 58 -39 63
rect -54 56 -39 58
rect -33 63 -18 65
rect -33 58 -28 63
rect -23 58 -18 63
rect -33 56 -18 58
rect -12 63 3 65
rect -12 58 -7 63
rect -2 58 3 63
rect -12 56 3 58
rect 9 63 24 65
rect 9 58 14 63
rect 19 58 24 63
rect 9 56 24 58
<< psubdiffcont >>
rect -49 -50 -44 -45
rect -28 -50 -23 -45
rect -7 -50 -2 -45
rect 14 -50 19 -45
<< nsubdiffcont >>
rect -49 58 -44 63
rect -28 58 -23 63
rect -7 58 -2 63
rect 14 58 19 63
<< polysilicon >>
rect -41 49 -35 54
rect -30 49 -24 54
rect -13 49 -7 54
rect 4 49 10 54
rect -41 3 -35 15
rect -45 1 -35 3
rect -45 -5 -43 1
rect -37 -5 -35 1
rect -45 -7 -35 -5
rect -30 3 -24 15
rect -13 3 -7 15
rect 4 3 10 15
rect -30 1 -19 3
rect -30 -5 -27 1
rect -21 -5 -19 1
rect -30 -7 -19 -5
rect -14 1 -3 3
rect -14 -5 -11 1
rect -5 -5 -3 1
rect -14 -7 -3 -5
rect 3 1 13 3
rect 3 -5 5 1
rect 11 -5 13 1
rect 3 -7 13 -5
rect -41 -19 -35 -7
rect -24 -14 -19 -7
rect -7 -10 -3 -7
rect -24 -19 -18 -14
rect -7 -19 -1 -10
rect 4 -19 10 -7
rect -41 -41 -35 -36
rect -24 -41 -18 -36
rect -7 -41 -1 -36
rect 4 -41 10 -36
<< polycontact >>
rect -43 -5 -37 1
rect -27 -5 -21 1
rect -11 -5 -5 1
rect 5 -5 11 1
<< metal1 >>
rect -60 63 29 70
rect -60 58 -49 63
rect -44 58 -28 63
rect -23 58 -7 63
rect -2 58 14 63
rect 19 58 29 63
rect -60 56 29 58
rect -49 47 -44 56
rect -49 37 -44 42
rect -4 47 1 56
rect -4 37 1 42
rect -49 30 -44 32
rect -21 34 -16 37
rect -4 30 1 32
rect 13 34 18 37
rect -21 24 -16 29
rect 13 24 18 29
rect -16 19 13 22
rect -21 17 18 19
rect 13 11 18 17
rect 13 6 26 11
rect 20 1 26 6
rect -45 -5 -43 1
rect -37 -5 -35 1
rect -29 -5 -27 1
rect -21 -5 -19 1
rect -13 -5 -11 1
rect -5 -5 -3 1
rect 3 -5 5 1
rect 11 -5 13 1
rect 19 0 27 1
rect 19 -6 20 0
rect 26 -6 27 0
rect 19 -7 27 -6
rect 20 -13 26 -7
rect -49 -19 -10 -14
rect -49 -23 -44 -19
rect -15 -23 -10 -19
rect -49 -33 -44 -31
rect -32 -26 -27 -24
rect -15 -33 -10 -31
rect 13 -19 26 -13
rect 13 -23 18 -19
rect 13 -33 18 -31
rect -32 -43 -27 -34
rect -60 -45 29 -43
rect -60 -50 -49 -45
rect -44 -50 -28 -45
rect -23 -50 -7 -45
rect -2 -50 14 -45
rect 19 -50 29 -45
rect -60 -57 29 -50
<< via1 >>
rect -43 -5 -37 1
rect -27 -5 -21 1
rect -11 -5 -5 1
rect 5 -5 11 1
rect 20 -6 26 0
<< metal2 >>
rect -45 1 -35 2
rect -45 -5 -43 1
rect -37 -5 -35 1
rect -45 -6 -35 -5
rect -29 1 -19 2
rect -29 -5 -27 1
rect -21 -5 -19 1
rect -29 -6 -19 -5
rect -13 1 -3 2
rect -13 -5 -11 1
rect -5 -5 -3 1
rect -13 -6 -3 -5
rect 3 1 13 2
rect 3 -5 5 1
rect 11 -5 13 1
rect 3 -6 13 -5
rect 19 0 27 1
rect 19 -6 20 0
rect 26 -6 27 0
rect 19 -7 27 -6
<< labels >>
rlabel via1 -40 -2 -40 -2 0 A0
rlabel metal2 -27 -5 -21 1 0 A1
rlabel metal2 -11 -5 -5 1 0 B
rlabel metal2 5 -5 11 1 0 C
rlabel metal2 20 -6 26 0 0 out
rlabel nsubdiffcont -49 58 -44 63 0 vdd
rlabel psubdiffcont -49 -50 -44 -45 0 vss
<< end >>
