magic
tech gf180mcuD
timestamp 1755140435
<< nwell >>
rect -6 44 106 122
<< nmos >>
rect 19 15 25 32
rect 30 15 36 32
rect 49 15 55 32
rect 68 15 74 32
rect 79 15 85 32
<< pmos >>
rect 13 68 19 102
rect 30 68 36 102
rect 47 68 53 102
rect 64 68 70 102
rect 81 68 87 102
<< ndiff >>
rect 9 29 19 32
rect 9 17 11 29
rect 16 17 19 29
rect 9 15 19 17
rect 25 15 30 32
rect 36 29 49 32
rect 36 17 39 29
rect 44 17 49 29
rect 36 15 49 17
rect 55 29 68 32
rect 55 17 60 29
rect 65 17 68 29
rect 55 15 68 17
rect 74 15 79 32
rect 85 29 95 32
rect 85 17 88 29
rect 93 17 95 29
rect 85 15 95 17
<< pdiff >>
rect 3 85 13 102
rect 3 80 5 85
rect 10 80 13 85
rect 3 75 13 80
rect 3 70 5 75
rect 10 70 13 75
rect 3 68 13 70
rect 19 98 30 102
rect 19 93 22 98
rect 27 93 30 98
rect 19 88 30 93
rect 19 83 22 88
rect 27 83 30 88
rect 19 68 30 83
rect 36 85 47 102
rect 36 80 39 85
rect 44 80 47 85
rect 36 75 47 80
rect 36 70 39 75
rect 44 70 47 75
rect 36 68 47 70
rect 53 99 64 102
rect 53 94 56 99
rect 61 94 64 99
rect 53 89 64 94
rect 53 84 56 89
rect 61 84 64 89
rect 53 68 64 84
rect 70 85 81 102
rect 70 80 73 85
rect 78 80 81 85
rect 70 75 81 80
rect 70 70 73 75
rect 78 70 81 75
rect 70 68 81 70
rect 87 99 97 102
rect 87 94 90 99
rect 95 94 97 99
rect 87 89 97 94
rect 87 84 90 89
rect 95 84 97 89
rect 87 68 97 84
<< ndiffc >>
rect 11 17 16 29
rect 39 17 44 29
rect 60 17 65 29
rect 88 17 93 29
<< pdiffc >>
rect 5 80 10 85
rect 5 70 10 75
rect 22 93 27 98
rect 22 83 27 88
rect 39 80 44 85
rect 39 70 44 75
rect 56 94 61 99
rect 56 84 61 89
rect 73 80 78 85
rect 73 70 78 75
rect 90 94 95 99
rect 90 84 95 89
<< psubdiff >>
rect 0 5 15 7
rect 0 0 4 5
rect 9 0 15 5
rect 0 -2 15 0
rect 21 5 36 7
rect 21 0 26 5
rect 31 0 36 5
rect 21 -2 36 0
rect 42 5 57 7
rect 42 0 47 5
rect 52 0 57 5
rect 42 -2 57 0
rect 63 5 78 7
rect 63 0 68 5
rect 73 0 78 5
rect 63 -2 78 0
rect 84 5 99 7
rect 84 0 89 5
rect 94 0 99 5
rect 84 -2 99 0
<< nsubdiff >>
rect 3 117 18 119
rect 3 112 8 117
rect 13 112 18 117
rect 3 110 18 112
rect 24 117 39 119
rect 24 112 29 117
rect 34 112 39 117
rect 24 110 39 112
rect 45 117 60 119
rect 45 112 50 117
rect 55 112 60 117
rect 45 110 60 112
rect 66 117 81 119
rect 66 112 71 117
rect 76 112 81 117
rect 66 110 81 112
<< psubdiffcont >>
rect 4 0 9 5
rect 26 0 31 5
rect 47 0 52 5
rect 68 0 73 5
rect 89 0 94 5
<< nsubdiffcont >>
rect 8 112 13 117
rect 29 112 34 117
rect 50 112 55 117
rect 71 112 76 117
<< polysilicon >>
rect 13 102 19 107
rect 30 102 36 107
rect 47 102 53 107
rect 64 102 70 107
rect 81 102 87 107
rect 13 63 19 68
rect 13 54 17 63
rect 6 50 17 54
rect 30 53 36 68
rect 47 54 53 68
rect 64 54 70 68
rect 81 63 87 68
rect 81 61 96 63
rect 81 60 97 61
rect 81 59 89 60
rect 86 55 89 59
rect 94 55 97 60
rect 25 51 36 53
rect 2 47 11 50
rect 2 42 4 47
rect 9 42 11 47
rect 25 46 29 51
rect 34 46 36 51
rect 25 44 36 46
rect 43 52 54 54
rect 43 47 47 52
rect 52 47 54 52
rect 43 45 54 47
rect 61 52 72 54
rect 86 53 97 55
rect 61 47 65 52
rect 70 47 72 52
rect 61 45 72 47
rect 2 40 11 42
rect 6 38 11 40
rect 6 34 25 38
rect 32 37 36 44
rect 19 32 25 34
rect 30 32 36 37
rect 49 37 53 45
rect 68 37 72 45
rect 81 49 96 53
rect 81 40 85 49
rect 49 32 55 37
rect 68 32 74 37
rect 79 32 85 40
rect 19 10 25 15
rect 30 10 36 15
rect 49 10 55 15
rect 68 10 74 15
rect 79 10 85 15
<< polycontact >>
rect 89 55 94 60
rect 4 42 9 47
rect 29 46 34 51
rect 47 47 52 52
rect 65 47 70 52
<< metal1 >>
rect -6 117 106 122
rect -6 112 8 117
rect 13 112 29 117
rect 34 112 50 117
rect 55 112 71 117
rect 76 112 106 117
rect -6 108 106 112
rect 22 98 27 108
rect 22 88 27 93
rect 5 85 10 87
rect 56 99 95 101
rect 61 96 90 99
rect 56 89 61 94
rect 22 80 27 83
rect 39 85 44 87
rect 90 89 95 94
rect 56 82 61 84
rect 73 85 78 87
rect 5 75 10 80
rect 5 63 10 70
rect 39 75 44 80
rect 39 63 44 70
rect 5 58 44 63
rect 90 82 95 84
rect 73 75 78 80
rect 73 62 78 70
rect 73 57 82 62
rect 2 48 11 49
rect -2 42 3 48
rect 9 42 11 48
rect 23 45 28 51
rect 34 45 36 51
rect 41 46 46 52
rect 52 46 54 52
rect 59 46 64 52
rect 70 46 72 52
rect 2 41 11 42
rect 77 41 82 57
rect 87 54 89 60
rect 95 54 97 60
rect 88 41 93 46
rect 39 36 93 41
rect 99 40 101 46
rect 11 29 16 31
rect 11 9 16 17
rect 39 29 44 36
rect 39 15 44 17
rect 60 29 65 31
rect 60 9 65 17
rect 88 29 93 36
rect 88 15 93 17
rect -6 5 106 9
rect -6 0 4 5
rect 9 0 26 5
rect 31 0 47 5
rect 52 0 68 5
rect 73 0 89 5
rect 94 0 106 5
rect -6 -5 106 0
<< via1 >>
rect 3 47 9 48
rect 3 42 4 47
rect 4 42 9 47
rect 28 46 29 51
rect 29 46 34 51
rect 28 45 34 46
rect 46 47 47 52
rect 47 47 52 52
rect 46 46 52 47
rect 64 47 65 52
rect 65 47 70 52
rect 64 46 70 47
rect 89 55 94 60
rect 94 55 95 60
rect 89 54 95 55
rect 93 40 99 46
<< metal2 >>
rect 87 60 97 61
rect 87 54 89 60
rect 95 54 97 60
rect 87 53 97 54
rect 43 52 54 53
rect 25 51 36 52
rect 0 48 11 49
rect 0 42 3 48
rect 9 42 11 48
rect 25 45 28 51
rect 34 45 36 51
rect 43 46 46 52
rect 52 46 54 52
rect 43 45 54 46
rect 61 52 72 53
rect 61 46 64 52
rect 70 46 72 52
rect 61 45 72 46
rect 90 46 101 47
rect 25 44 36 45
rect 0 41 11 42
rect 90 40 93 46
rect 99 40 101 46
rect 90 39 101 40
<< labels >>
rlabel metal1 -6 114 -6 114 3 vdd
rlabel metal1 -6 1 -6 1 3 vss
rlabel polysilicon 36 40 36 40 1 B0
rlabel polysilicon 68 42 68 42 1 A1
rlabel polysilicon 49 42 49 42 1 C
rlabel polysilicon 2 40 2 40 1 B1
rlabel polysilicon 85 42 85 42 1 A0
rlabel via1 95 40 95 40 1 Y
<< end >>
