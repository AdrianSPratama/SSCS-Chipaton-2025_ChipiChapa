* SPICE3 file created from gf180mcu_gp9t3v3__aoi221_1.ext - technology: gf180mcuD

X0 a_30_670# B0 vdd vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1 Y A1 a_530_670# vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X2 a_250_160# B1 vss vss nfet_03v3 ad=0.10625p pd=1.1u as=0.425p ps=2.7u w=0.85u l=0.3u
X3 vss C Y vss nfet_03v3 ad=0.27625p pd=1.5u as=0.27625p ps=1.5u w=0.85u l=0.3u
X4 a_530_670# A0 Y vdd pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X5 Y A0 a_740_160# vss nfet_03v3 ad=0.425p pd=2.7u as=0.10625p ps=1.1u w=0.85u l=0.3u
X6 vdd B1 a_30_670# vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.85p ps=4.4u w=1.7u l=0.3u
X7 Y B0 a_250_160# vss nfet_03v3 ad=0.27625p pd=1.5u as=0.10625p ps=1.1u w=0.85u l=0.3u
X8 a_740_160# A1 vss vss nfet_03v3 ad=0.10625p pd=1.1u as=0.27625p ps=1.5u w=0.85u l=0.3u
X9 a_530_670# C a_30_670# vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
C0 a_530_670# A1 0.03341f
C1 C Y 0.13459f
C2 C vdd 0.10597f
C3 A0 a_530_670# 0.04623f
C4 Y B1 0.00897f
C5 vdd B1 0.10787f
C6 A1 Y 0.21331f
C7 vdd A1 0.08965f
C8 A0 vdd 0.12702f
C9 A0 Y 0.21193f
C10 B0 a_30_670# 0.1005f
C11 a_530_670# a_30_670# 0.02429f
C12 a_530_670# B0 0.00134f
C13 a_30_670# Y 0.04804f
C14 vdd a_30_670# 0.17787f
C15 B0 Y 0.00974f
C16 B0 vdd 0.10252f
C17 C B1 0
C18 a_530_670# Y 0.10318f
C19 a_530_670# vdd 0.26686f
C20 C A1 0.11332f
C21 A0 C 0
C22 A1 B1 0
C23 A0 B1 0
C24 vdd Y 0.02607f
C25 A0 A1 0.07085f
C26 a_30_670# a_250_160# 0
C27 B0 a_250_160# 0.00221f
C28 C a_30_670# 0.01213f
C29 a_30_670# B1 0.08494f
C30 B0 C 0.10697f
C31 a_30_670# A1 0.00307f
C32 Y a_740_160# 0.0043f
C33 A0 a_30_670# 0
C34 B0 B1 0.11641f
C35 Y a_250_160# 0
C36 a_530_670# C 0.00502f
C37 B0 A1 0
C38 A0 B0 0
C39 Y vss 0.57547f
C40 A0 vss 0.37725f
C41 A1 vss 0.29923f
C42 C vss 0.29661f
C43 B0 vss 0.30231f
C44 B1 vss 0.43242f
C45 vdd vss 2.41757f
C46 a_740_160# vss 0.00366f
C47 a_250_160# vss 0.00366f
C48 a_530_670# vss 0.05393f
C49 a_30_670# vss 0.09822f
