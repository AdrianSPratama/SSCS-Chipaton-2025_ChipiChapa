VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp9t3v3_aoi211_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3_aoi211_1 ;
  ORIGIN 0.900 0.900 ;
  SIZE 4.450 BY 6.350 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -0.900 2.250 3.550 5.450 ;
      LAYER Metal1 ;
        RECT -0.900 4.750 3.550 5.450 ;
        RECT 0.500 3.300 0.750 4.750 ;
    END
  END vdd
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 1.750 1.200 2.050 ;
      LAYER Metal2 ;
        RECT 0.700 1.700 1.200 2.100 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT -0.150 1.750 0.350 2.050 ;
      LAYER Metal2 ;
        RECT -0.150 1.700 0.350 2.100 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.500 1.750 2.000 2.050 ;
      LAYER Metal2 ;
        RECT 1.500 1.700 2.000 2.100 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.765000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.300 1.750 2.800 2.050 ;
      LAYER Metal2 ;
        RECT 2.300 1.700 2.800 2.100 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.742500 ;
    PORT
      LAYER Metal1 ;
        RECT 2.750 2.600 3.000 3.700 ;
        RECT 2.750 2.300 3.300 2.600 ;
        RECT 3.050 2.100 3.300 2.300 ;
        RECT 3.050 1.700 3.550 2.100 ;
        RECT 3.050 1.400 3.300 1.700 ;
        RECT 1.350 1.150 3.300 1.400 ;
        RECT 1.350 0.250 1.600 1.150 ;
        RECT 3.050 0.250 3.300 1.150 ;
      LAYER Metal2 ;
        RECT 3.150 1.700 3.550 2.100 ;
    END
  END Y
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT -0.350 -0.200 -0.100 0.900 ;
        RECT 2.200 -0.200 2.450 0.900 ;
        RECT -0.900 -0.900 3.550 -0.200 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT -0.350 3.000 -0.100 3.950 ;
        RECT 1.350 3.000 1.600 3.950 ;
        RECT -0.350 2.750 1.600 3.000 ;
  END
END gf180mcu_osu_sc_gp9t3v3_aoi211_1
END LIBRARY

