magic
tech gf180mcuD
timestamp 1758084589
<< nwell >>
rect -6 58 106 122
<< nmos >>
rect 17 16 23 33
rect 30 16 36 33
rect 47 16 53 33
rect 64 16 70 33
rect 77 16 83 33
<< pmos >>
rect 13 67 19 101
rect 30 67 36 101
rect 47 67 53 101
rect 64 67 70 101
rect 81 67 87 101
<< ndiff >>
rect 7 31 17 33
rect 7 18 9 31
rect 14 18 17 31
rect 7 16 17 18
rect 23 16 30 33
rect 36 31 47 33
rect 36 18 39 31
rect 44 18 47 31
rect 36 16 47 18
rect 53 31 64 33
rect 53 18 56 31
rect 61 18 64 31
rect 53 16 64 18
rect 70 16 77 33
rect 83 31 93 33
rect 83 18 86 31
rect 91 18 93 31
rect 83 16 93 18
<< pdiff >>
rect 3 99 13 101
rect 3 74 5 99
rect 10 74 13 99
rect 3 67 13 74
rect 19 99 30 101
rect 19 79 22 99
rect 27 79 30 99
rect 19 67 30 79
rect 36 99 47 101
rect 36 74 39 99
rect 44 74 47 99
rect 36 67 47 74
rect 53 94 64 101
rect 53 69 56 94
rect 61 69 64 94
rect 53 67 64 69
rect 70 89 81 101
rect 70 75 73 89
rect 78 75 81 89
rect 70 67 81 75
rect 87 94 97 101
rect 87 80 90 94
rect 95 80 97 94
rect 87 67 97 80
<< ndiffc >>
rect 9 18 14 31
rect 39 18 44 31
rect 56 18 61 31
rect 86 18 91 31
<< pdiffc >>
rect 5 74 10 99
rect 22 79 27 99
rect 39 74 44 99
rect 56 69 61 94
rect 73 75 78 89
rect 90 80 95 94
<< psubdiff >>
rect 0 7 15 9
rect 0 2 5 7
rect 10 2 15 7
rect 0 0 15 2
rect 21 7 36 9
rect 21 2 26 7
rect 31 2 36 7
rect 21 0 36 2
rect 42 7 57 9
rect 42 2 47 7
rect 52 2 57 7
rect 42 0 57 2
rect 63 7 78 9
rect 63 2 68 7
rect 73 2 78 7
rect 63 0 78 2
rect 84 7 99 9
rect 84 2 89 7
rect 94 2 99 7
rect 84 0 99 2
<< nsubdiff >>
rect 0 115 15 117
rect 0 110 5 115
rect 10 110 15 115
rect 0 108 15 110
rect 21 115 36 117
rect 21 110 26 115
rect 31 110 36 115
rect 21 108 36 110
rect 42 115 57 117
rect 42 110 47 115
rect 52 110 57 115
rect 42 108 57 110
rect 63 115 78 117
rect 63 110 68 115
rect 73 110 78 115
rect 63 108 78 110
rect 84 115 99 117
rect 84 110 89 115
rect 94 110 99 115
rect 84 108 99 110
<< psubdiffcont >>
rect 5 2 10 7
rect 26 2 31 7
rect 47 2 52 7
rect 68 2 73 7
rect 89 2 94 7
<< nsubdiffcont >>
rect 5 110 10 115
rect 26 110 31 115
rect 47 110 52 115
rect 68 110 73 115
rect 89 110 94 115
<< polysilicon >>
rect 13 101 19 106
rect 30 101 36 106
rect 47 101 53 106
rect 64 101 70 106
rect 81 101 87 106
rect 13 62 19 67
rect 30 62 36 67
rect 47 62 53 67
rect 64 62 70 67
rect 81 62 87 67
rect 13 60 23 62
rect 13 54 15 60
rect 21 54 23 60
rect 13 52 23 54
rect 29 60 39 62
rect 29 54 31 60
rect 37 54 39 60
rect 29 52 39 54
rect 45 60 55 62
rect 45 54 47 60
rect 53 54 55 60
rect 45 52 55 54
rect 61 60 71 62
rect 61 54 63 60
rect 69 54 71 60
rect 61 52 71 54
rect 77 60 87 62
rect 77 54 79 60
rect 85 54 87 60
rect 77 52 87 54
rect 17 33 23 52
rect 30 33 36 52
rect 47 33 53 52
rect 64 33 70 52
rect 77 33 83 52
rect 17 11 23 16
rect 30 11 36 16
rect 47 11 53 16
rect 64 11 70 16
rect 77 11 83 16
<< polycontact >>
rect 15 54 21 60
rect 31 54 37 60
rect 47 54 53 60
rect 63 54 69 60
rect 79 54 85 60
<< metal1 >>
rect -6 115 106 122
rect -6 110 5 115
rect 10 110 26 115
rect 31 110 47 115
rect 52 110 68 115
rect 73 110 89 115
rect 94 110 106 115
rect -6 108 106 110
rect 5 99 10 101
rect 22 99 27 108
rect 22 77 27 79
rect 39 99 44 101
rect 5 72 10 74
rect 39 72 44 74
rect 5 67 44 72
rect 56 96 95 101
rect 56 94 61 96
rect 90 94 95 96
rect 56 67 61 69
rect 73 89 78 91
rect 90 78 95 80
rect 73 73 78 75
rect 73 67 98 73
rect 13 54 15 60
rect 21 54 23 60
rect 29 54 31 60
rect 37 54 39 60
rect 45 54 47 60
rect 53 54 55 60
rect 61 54 63 60
rect 69 54 71 60
rect 77 54 79 60
rect 85 54 87 60
rect 92 47 98 67
rect 39 41 92 47
rect 98 41 100 47
rect 9 31 14 33
rect 9 9 14 18
rect 39 31 44 41
rect 39 16 44 18
rect 56 31 61 33
rect 56 9 61 18
rect 86 31 91 41
rect 86 16 91 18
rect -6 7 106 9
rect -6 2 5 7
rect 10 2 26 7
rect 31 2 47 7
rect 52 2 68 7
rect 73 2 89 7
rect 94 2 106 7
rect -6 -5 106 2
<< via1 >>
rect 15 54 21 60
rect 31 54 37 60
rect 47 54 53 60
rect 63 54 69 60
rect 79 54 85 60
rect 92 41 98 47
<< metal2 >>
rect 13 60 23 61
rect 13 54 15 60
rect 21 54 23 60
rect 13 53 23 54
rect 29 60 39 61
rect 29 54 31 60
rect 37 54 39 60
rect 29 53 39 54
rect 45 60 55 61
rect 45 54 47 60
rect 53 54 55 60
rect 45 53 55 54
rect 61 60 71 61
rect 61 54 63 60
rect 69 54 71 60
rect 61 53 71 54
rect 77 60 87 61
rect 77 54 79 60
rect 85 54 87 60
rect 77 53 87 54
rect 91 47 99 48
rect 91 41 92 47
rect 98 41 99 47
rect 91 40 99 41
<< labels >>
rlabel metal1 -6 114 -6 114 3 vdd
port 7 e power bidirectional abutment
rlabel metal1 -6 1 -6 1 3 vss
port 8 e ground bidirectional abutment
rlabel polycontact 82 57 82 57 1 A0
port 1 n signal input
rlabel via1 94 41 94 41 1 Y
port 6 n signal output
rlabel polycontact 66 57 66 57 1 A1
port 2 n signal input
rlabel polycontact 50 57 50 57 1 C
port 5 n signal input
rlabel polycontact 34 57 34 57 1 B0
port 3 n signal input
rlabel polycontact 18 57 18 57 1 B1
port 4 n signal input
<< end >>
