magic
tech gf180mcuD
timestamp 1757698147
<< nwell >>
rect -60 4 29 68
<< nmos >>
rect -41 -38 -35 -21
rect -24 -38 -18 -21
rect -7 -38 -1 -21
rect 4 -38 10 -21
<< pmos >>
rect -41 13 -35 47
rect -30 13 -24 47
rect -13 13 -7 47
rect 4 13 10 47
<< ndiff >>
rect -51 -25 -41 -21
rect -51 -33 -49 -25
rect -44 -33 -41 -25
rect -51 -38 -41 -33
rect -35 -28 -24 -21
rect -35 -36 -32 -28
rect -27 -36 -24 -28
rect -35 -38 -24 -36
rect -18 -25 -7 -21
rect -18 -33 -15 -25
rect -10 -33 -7 -25
rect -18 -38 -7 -33
rect -1 -38 4 -21
rect 10 -25 20 -21
rect 10 -33 13 -25
rect 18 -33 20 -25
rect 10 -38 20 -33
<< pdiff >>
rect -51 45 -41 47
rect -51 40 -49 45
rect -44 40 -41 45
rect -51 35 -41 40
rect -51 30 -49 35
rect -44 30 -41 35
rect -51 13 -41 30
rect -35 13 -30 47
rect -24 32 -13 47
rect -24 27 -21 32
rect -16 27 -13 32
rect -24 22 -13 27
rect -24 17 -21 22
rect -16 17 -13 22
rect -24 13 -13 17
rect -7 45 4 47
rect -7 40 -4 45
rect 1 40 4 45
rect -7 35 4 40
rect -7 30 -4 35
rect 1 30 4 35
rect -7 13 4 30
rect 10 32 20 47
rect 10 27 13 32
rect 18 27 20 32
rect 10 22 20 27
rect 10 17 13 22
rect 18 17 20 22
rect 10 13 20 17
<< ndiffc >>
rect -49 -33 -44 -25
rect -32 -36 -27 -28
rect -15 -33 -10 -25
rect 13 -33 18 -25
<< pdiffc >>
rect -49 40 -44 45
rect -49 30 -44 35
rect -21 27 -16 32
rect -21 17 -16 22
rect -4 40 1 45
rect -4 30 1 35
rect 13 27 18 32
rect 13 17 18 22
<< psubdiff >>
rect -54 -47 -39 -45
rect -54 -52 -49 -47
rect -44 -52 -39 -47
rect -54 -54 -39 -52
rect -33 -47 -18 -45
rect -33 -52 -28 -47
rect -23 -52 -18 -47
rect -33 -54 -18 -52
rect -12 -47 3 -45
rect -12 -52 -7 -47
rect -2 -52 3 -47
rect -12 -54 3 -52
rect 9 -47 24 -45
rect 9 -52 14 -47
rect 19 -52 24 -47
rect 9 -54 24 -52
<< nsubdiff >>
rect -54 61 -39 63
rect -54 56 -49 61
rect -44 56 -39 61
rect -54 54 -39 56
rect -33 61 -18 63
rect -33 56 -28 61
rect -23 56 -18 61
rect -33 54 -18 56
rect -12 61 3 63
rect -12 56 -7 61
rect -2 56 3 61
rect -12 54 3 56
rect 9 61 24 63
rect 9 56 14 61
rect 19 56 24 61
rect 9 54 24 56
<< psubdiffcont >>
rect -49 -52 -44 -47
rect -28 -52 -23 -47
rect -7 -52 -2 -47
rect 14 -52 19 -47
<< nsubdiffcont >>
rect -49 56 -44 61
rect -28 56 -23 61
rect -7 56 -2 61
rect 14 56 19 61
<< polysilicon >>
rect -41 47 -35 52
rect -30 47 -24 52
rect -13 47 -7 52
rect 4 47 10 52
rect -41 11 -35 13
rect -46 8 -35 11
rect -52 7 -35 8
rect -30 8 -24 13
rect -13 8 -7 13
rect 4 8 10 13
rect -52 6 -42 7
rect -52 0 -50 6
rect -44 0 -42 6
rect -52 -2 -42 0
rect -46 -12 -42 -2
rect -30 6 -20 8
rect -30 0 -28 6
rect -22 0 -20 6
rect -30 -2 -20 0
rect -14 6 -4 8
rect -14 0 -12 6
rect -6 0 -4 6
rect -14 -2 -4 0
rect 2 6 12 8
rect 2 0 4 6
rect 10 0 12 6
rect 2 -2 12 0
rect -30 -12 -24 -2
rect -12 -12 -7 -2
rect -46 -16 -35 -12
rect -30 -16 -20 -12
rect -12 -16 -1 -12
rect -41 -21 -35 -16
rect -24 -21 -18 -16
rect -7 -21 -1 -16
rect 4 -21 10 -2
rect -41 -43 -35 -38
rect -24 -43 -18 -38
rect -7 -43 -1 -38
rect 4 -43 10 -38
<< polycontact >>
rect -50 0 -44 6
rect -28 0 -22 6
rect -12 0 -6 6
rect 4 0 10 6
<< metal1 >>
rect -60 61 29 68
rect -60 56 -49 61
rect -44 56 -28 61
rect -23 56 -7 61
rect -2 56 14 61
rect 19 56 29 61
rect -60 54 29 56
rect -49 45 -44 54
rect -49 35 -44 40
rect -4 45 1 54
rect -4 35 1 40
rect -49 28 -44 30
rect -21 32 -16 35
rect -4 28 1 30
rect 13 32 18 35
rect -21 22 -16 27
rect 13 22 18 27
rect -16 17 13 20
rect -21 16 18 17
rect -21 15 24 16
rect 13 11 24 15
rect -52 0 -50 6
rect -44 0 -42 6
rect -30 0 -28 6
rect -22 0 -20 6
rect -14 0 -12 6
rect -6 0 -4 6
rect 2 0 4 6
rect 10 0 12 6
rect 19 -6 24 11
rect 16 -7 24 -6
rect 16 -13 17 -7
rect 23 -13 24 -7
rect 16 -14 24 -13
rect -49 -21 -10 -16
rect -49 -25 -44 -21
rect -15 -25 -10 -21
rect -49 -35 -44 -33
rect -32 -28 -27 -26
rect -15 -35 -10 -33
rect 13 -19 24 -14
rect 13 -25 18 -19
rect 13 -35 18 -33
rect -32 -45 -27 -36
rect -60 -47 29 -45
rect -60 -52 -49 -47
rect -44 -52 -28 -47
rect -23 -52 -7 -47
rect -2 -52 14 -47
rect 19 -52 29 -47
rect -60 -59 29 -52
<< via1 >>
rect -50 0 -44 6
rect -28 0 -22 6
rect -12 0 -6 6
rect 4 0 10 6
rect 17 -13 23 -7
<< metal2 >>
rect -52 6 -42 7
rect -52 0 -50 6
rect -44 0 -42 6
rect -52 -1 -42 0
rect -30 6 -20 7
rect -30 0 -28 6
rect -22 0 -20 6
rect -30 -1 -20 0
rect -14 6 -4 7
rect -14 0 -12 6
rect -6 0 -4 6
rect -14 -1 -4 0
rect 2 6 12 7
rect 2 0 4 6
rect 10 0 12 6
rect 2 -1 12 0
rect 16 -7 24 -6
rect 16 -13 17 -7
rect 23 -13 24 -7
rect 16 -14 24 -13
<< labels >>
rlabel nsubdiffcont -49 56 -44 61 0 vdd
port 6 n power bidirectional abutment
rlabel psubdiffcont -49 -52 -44 -47 0 vss
port 7 s ground bidirectional abutment
rlabel metal2 -50 0 -44 6 0 A0
port 1 w signal input
rlabel metal2 17 -13 23 -7 0 Y
port 5 e signal output
rlabel metal2 4 0 10 6 0 C
port 4 w signal input
rlabel metal2 -12 0 -6 6 0 B
port 3 w signal input
rlabel metal2 -28 0 -22 6 0 A1
port 2 w signal input
<< end >>
