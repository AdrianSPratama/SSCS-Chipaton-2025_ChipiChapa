magic
tech gf180mcuD
timestamp 1757661659
<< nwell >>
rect -60 6 29 70
<< nmos >>
rect -41 -36 -35 -19
rect -24 -36 -18 -19
rect -7 -36 -1 -19
rect 4 -36 10 -19
<< pmos >>
rect -41 15 -35 49
rect -30 15 -24 49
rect -13 15 -7 49
rect 4 15 10 49
<< ndiff >>
rect -51 -23 -41 -19
rect -51 -31 -49 -23
rect -44 -31 -41 -23
rect -51 -36 -41 -31
rect -35 -26 -24 -19
rect -35 -34 -32 -26
rect -27 -34 -24 -26
rect -35 -36 -24 -34
rect -18 -23 -7 -19
rect -18 -31 -15 -23
rect -10 -31 -7 -23
rect -18 -36 -7 -31
rect -1 -36 4 -19
rect 10 -23 20 -19
rect 10 -31 13 -23
rect 18 -31 20 -23
rect 10 -36 20 -31
<< pdiff >>
rect -51 47 -41 49
rect -51 42 -49 47
rect -44 42 -41 47
rect -51 37 -41 42
rect -51 32 -49 37
rect -44 32 -41 37
rect -51 15 -41 32
rect -35 15 -30 49
rect -24 34 -13 49
rect -24 29 -21 34
rect -16 29 -13 34
rect -24 24 -13 29
rect -24 19 -21 24
rect -16 19 -13 24
rect -24 15 -13 19
rect -7 47 4 49
rect -7 42 -4 47
rect 1 42 4 47
rect -7 37 4 42
rect -7 32 -4 37
rect 1 32 4 37
rect -7 15 4 32
rect 10 34 20 49
rect 10 29 13 34
rect 18 29 20 34
rect 10 24 20 29
rect 10 19 13 24
rect 18 19 20 24
rect 10 15 20 19
<< ndiffc >>
rect -49 -31 -44 -23
rect -32 -34 -27 -26
rect -15 -31 -10 -23
rect 13 -31 18 -23
<< pdiffc >>
rect -49 42 -44 47
rect -49 32 -44 37
rect -21 29 -16 34
rect -21 19 -16 24
rect -4 42 1 47
rect -4 32 1 37
rect 13 29 18 34
rect 13 19 18 24
<< psubdiff >>
rect -54 -45 -39 -43
rect -54 -50 -49 -45
rect -44 -50 -39 -45
rect -54 -52 -39 -50
rect -33 -45 -18 -43
rect -33 -50 -28 -45
rect -23 -50 -18 -45
rect -33 -52 -18 -50
rect -12 -45 3 -43
rect -12 -50 -7 -45
rect -2 -50 3 -45
rect -12 -52 3 -50
rect 9 -45 24 -43
rect 9 -50 14 -45
rect 19 -50 24 -45
rect 9 -52 24 -50
<< nsubdiff >>
rect -54 63 -39 65
rect -54 58 -49 63
rect -44 58 -39 63
rect -54 56 -39 58
rect -33 63 -18 65
rect -33 58 -28 63
rect -23 58 -18 63
rect -33 56 -18 58
rect -12 63 3 65
rect -12 58 -7 63
rect -2 58 3 63
rect -12 56 3 58
rect 9 63 24 65
rect 9 58 14 63
rect 19 58 24 63
rect 9 56 24 58
<< psubdiffcont >>
rect -49 -50 -44 -45
rect -28 -50 -23 -45
rect -7 -50 -2 -45
rect 14 -50 19 -45
<< nsubdiffcont >>
rect -49 58 -44 63
rect -28 58 -23 63
rect -7 58 -2 63
rect 14 58 19 63
<< polysilicon >>
rect -41 49 -35 54
rect -30 49 -24 54
rect -13 49 -7 54
rect 4 49 10 54
rect -41 13 -35 15
rect -46 9 -35 13
rect -46 8 -42 9
rect -52 6 -42 8
rect -52 0 -50 6
rect -44 0 -42 6
rect -52 -2 -42 0
rect -46 -10 -42 -2
rect -30 8 -24 15
rect -13 8 -7 15
rect 4 8 10 15
rect -30 6 -20 8
rect -30 0 -28 6
rect -22 0 -20 6
rect -30 -2 -20 0
rect -14 6 -4 8
rect -14 0 -12 6
rect -6 0 -4 6
rect -14 -2 -4 0
rect 2 6 12 8
rect 2 0 4 6
rect 10 0 12 6
rect 2 -2 12 0
rect -30 -10 -24 -2
rect -12 -10 -7 -2
rect -46 -14 -35 -10
rect -30 -14 -20 -10
rect -12 -14 -1 -10
rect -41 -19 -35 -14
rect -24 -19 -18 -14
rect -7 -19 -1 -14
rect 4 -19 10 -2
rect -41 -41 -35 -36
rect -24 -41 -18 -36
rect -7 -41 -1 -36
rect 4 -41 10 -36
<< polycontact >>
rect -50 0 -44 6
rect -28 0 -22 6
rect -12 0 -6 6
rect 4 0 10 6
<< metal1 >>
rect -60 63 29 70
rect -60 58 -49 63
rect -44 58 -28 63
rect -23 58 -7 63
rect -2 58 14 63
rect 19 58 29 63
rect -60 56 29 58
rect -49 47 -44 56
rect -49 37 -44 42
rect -4 47 1 56
rect -4 37 1 42
rect -49 30 -44 32
rect -21 34 -16 37
rect -4 30 1 32
rect 13 34 18 37
rect -21 24 -16 29
rect 13 24 18 29
rect -16 19 13 22
rect -21 17 18 19
rect 13 16 18 17
rect 13 11 24 16
rect -52 0 -50 6
rect -44 0 -42 6
rect -30 0 -28 6
rect -22 0 -20 6
rect -14 0 -12 6
rect -6 0 -4 6
rect 2 0 4 6
rect 10 0 12 6
rect 19 -6 24 11
rect 16 -7 24 -6
rect 16 -13 17 -7
rect 23 -13 24 -7
rect -49 -19 -10 -14
rect -49 -23 -44 -19
rect -15 -23 -10 -19
rect -49 -33 -44 -31
rect -32 -26 -27 -24
rect -15 -33 -10 -31
rect 13 -19 24 -13
rect 13 -23 18 -19
rect 13 -33 18 -31
rect -32 -43 -27 -34
rect -60 -45 29 -43
rect -60 -50 -49 -45
rect -44 -50 -28 -45
rect -23 -50 -7 -45
rect -2 -50 14 -45
rect 19 -50 29 -45
rect -60 -57 29 -50
<< via1 >>
rect -50 0 -44 6
rect -28 0 -22 6
rect -12 0 -6 6
rect 4 0 10 6
rect 17 -13 23 -7
<< metal2 >>
rect -52 6 -42 7
rect -52 0 -50 6
rect -44 0 -42 6
rect -52 -1 -42 0
rect -30 6 -20 7
rect -30 0 -28 6
rect -22 0 -20 6
rect -30 -1 -20 0
rect -14 6 -4 7
rect -14 0 -12 6
rect -6 0 -4 6
rect -14 -1 -4 0
rect 2 6 12 7
rect 2 0 4 6
rect 10 0 12 6
rect 2 -1 12 0
rect 16 -7 24 -6
rect 16 -13 17 -7
rect 23 -13 24 -7
rect 16 -14 24 -13
<< labels >>
rlabel nsubdiffcont -49 58 -44 63 0 vdd
port 6 n power bidirectional abutment
rlabel psubdiffcont -49 -50 -44 -45 0 vss
port 7 s ground bidirectional abutment
rlabel metal2 17 -13 23 -7 0 Y
port 5 e signal output
rlabel metal2 4 0 10 6 0 C
port 4 w signal input
rlabel metal2 -12 0 -6 6 0 B
port 3 w signal input
rlabel metal2 -28 0 -22 6 0 A1
port 2 w signal input
rlabel metal2 -50 0 -44 6 0 A0
port 1 w signal input
<< end >>
