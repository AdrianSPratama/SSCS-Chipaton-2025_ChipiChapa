magic
tech gf180mcuD
timestamp 1755224193
use gf180mcu_gp9t3v3__aoi221_1  gf180mcu_gp9t3v3__aoi221_1_0
timestamp 1755140435
transform 1 0 107 0 1 5
box -6 -5 106 122
use gf180mcu_gp9t3v3_oai211_1  gf180mcu_gp9t3v3_oai211_1_0 /foss/designs/SSCS-Chipaton-2025_ChipiChapa/designs/oai211
timestamp 1755145353
transform 1 0 285 0 1 57
box -60 -57 29 70
use gf180mcu_gp9t3v3_oai221_1  gf180mcu_gp9t3v3_oai221_1_0 /foss/designs/SSCS-Chipaton-2025_ChipiChapa/designs/oai221
timestamp 1755166701
transform 1 0 343 0 1 31
box -17 -31 88 96
use gf180mcu_osu_sc_gp9t3v3_aoi211_1  gf180mcu_osu_sc_gp9t3v3_aoi211_1_0 /foss/designs/SSCS-Chipaton-2025_ChipiChapa/designs/aoi211
timestamp 1755166654
transform 1 0 18 0 1 18
box -18 -18 71 109
<< end >>
