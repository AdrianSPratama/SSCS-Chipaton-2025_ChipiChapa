* NGSPICE file created from gf180mcu_gp9t3v3_oai211_1.ext - technology: gf180mcuD

.subckt gf180mcu_gp9t3v3_oai211_1 A0 A1 B C Y vdd vss
X0 Y C vdd vdd pfet_03v3 ad=0.85p pd=4.4u as=0.4675p ps=2.25u w=1.7u l=0.3u
X1 a_n350_150# A0 vdd vdd pfet_03v3 ad=0.2125p pd=1.95u as=0.85p ps=4.4u w=1.7u l=0.3u
X2 a_n510_n360# A1 vss vss nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3 Y C a_n10_n360# vss nfet_03v3 ad=0.425p pd=2.7u as=0.10625p ps=1.1u w=0.85u l=0.3u
X4 Y A1 a_n350_150# vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.2125p ps=1.95u w=1.7u l=0.3u
X5 vdd B Y vdd pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X6 vss A0 a_n510_n360# vss nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X7 a_n10_n360# B a_n510_n360# vss nfet_03v3 ad=0.10625p pd=1.1u as=0.23375p ps=1.4u w=0.85u l=0.3u
C0 a_n350_150# a_n510_n360# 0.00253f
C1 A0 vdd 0.15557f
C2 C Y 0.1348f
C3 B vdd 0.10815f
C4 A0 A1 0.11598f
C5 A0 a_n510_n360# 0.05694f
C6 B A1 0.14363f
C7 B a_n510_n360# 0.02529f
C8 B C 0.16584f
C9 a_n10_n360# a_n510_n360# 0.00112f
C10 A1 vdd 0.10679f
C11 vdd a_n510_n360# 0.01096f
C12 a_n350_150# Y 0.00202f
C13 A1 a_n510_n360# 0.0593f
C14 a_n10_n360# C 0.00139f
C15 vdd C 0.11068f
C16 A0 Y 0.00474f
C17 B Y 0.07819f
C18 C a_n510_n360# 0.00287f
C19 a_n10_n360# Y 0.00189f
C20 vdd Y 0.23345f
C21 A1 Y 0.01598f
C22 a_n510_n360# Y 0.04443f
C23 a_n350_150# vdd 0.00727f
C24 Y vss 0.31065f
C25 C vss 0.33699f
C26 B vss 0.29561f
C27 A1 vss 0.30596f
C28 A0 vss 0.39977f
C29 vdd vss 1.96156f
C30 a_n10_n360# vss 0.00315f
C31 a_n510_n360# vss 0.3042f
.ends

