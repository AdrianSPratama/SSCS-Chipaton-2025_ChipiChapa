magic
tech gf180mcuC
timestamp 1753240757
<< nwell >>
rect 0 41 100 122
<< nmos >>
rect 12 12 18 32
rect 23 12 29 32
rect 40 12 46 32
rect 51 12 57 32
rect 70 17 76 27
<< pmos >>
rect 19 60 25 105
rect 36 60 42 105
rect 53 60 59 105
rect 70 60 76 105
<< ndiff >>
rect 2 28 12 32
rect 2 16 4 28
rect 9 16 12 28
rect 2 12 12 16
rect 18 12 23 32
rect 29 28 40 32
rect 29 16 32 28
rect 37 16 40 28
rect 29 12 40 16
rect 46 12 51 32
rect 57 28 68 32
rect 57 16 60 28
rect 65 27 68 28
rect 65 17 70 27
rect 76 25 86 27
rect 76 19 79 25
rect 84 19 86 25
rect 76 17 86 19
rect 65 16 68 17
rect 57 12 68 16
<< pdiff >>
rect 9 78 19 105
rect 9 73 11 78
rect 16 73 19 78
rect 9 68 19 73
rect 9 63 11 68
rect 16 63 19 68
rect 9 60 19 63
rect 25 101 36 105
rect 25 96 28 101
rect 33 96 36 101
rect 25 91 36 96
rect 25 86 28 91
rect 33 86 36 91
rect 25 60 36 86
rect 42 78 53 105
rect 42 73 45 78
rect 50 73 53 78
rect 42 68 53 73
rect 42 63 45 68
rect 50 63 53 68
rect 42 60 53 63
rect 59 60 70 105
rect 76 78 86 105
rect 76 73 79 78
rect 84 73 86 78
rect 76 68 86 73
rect 76 63 79 68
rect 84 63 86 68
rect 76 60 86 63
<< ndiffc >>
rect 4 16 9 28
rect 32 16 37 28
rect 60 16 65 28
rect 79 19 84 25
<< pdiffc >>
rect 11 73 16 78
rect 11 63 16 68
rect 28 96 33 101
rect 28 86 33 91
rect 45 73 50 78
rect 45 63 50 68
rect 79 73 84 78
rect 79 63 84 68
<< polysilicon >>
rect 19 105 25 110
rect 36 105 42 110
rect 53 105 59 110
rect 70 105 76 110
rect 19 55 25 60
rect 36 55 42 60
rect 53 55 59 60
rect 70 55 76 60
rect 12 32 18 37
rect 23 32 29 37
rect 40 32 46 37
rect 51 32 57 37
rect 72 32 76 37
rect 70 27 76 32
rect 70 12 76 17
rect 12 7 18 12
rect 23 7 29 12
rect 40 7 46 12
rect 51 7 57 12
<< metal1 >>
rect 0 108 100 122
rect 28 101 33 108
rect 28 91 33 96
rect 28 83 33 86
rect 11 78 16 80
rect 11 68 16 73
rect 11 62 16 63
rect 45 78 50 80
rect 45 68 50 73
rect 45 62 50 63
rect 79 78 84 80
rect 79 68 84 73
rect 79 62 84 63
rect 11 57 84 62
rect 32 35 84 40
rect 4 28 9 30
rect 4 9 9 16
rect 32 28 37 35
rect 32 14 37 16
rect 60 28 65 30
rect 79 25 84 35
rect 79 17 84 19
rect 60 9 65 16
rect 0 -5 100 9
<< labels >>
rlabel metal1 0 113 0 113 3 vdd
rlabel metal1 0 2 0 2 3 vss
rlabel polysilicon 12 33 12 33 1 A2
rlabel polysilicon 23 33 23 33 1 A1
rlabel polysilicon 40 33 40 33 1 B1
rlabel polysilicon 51 33 51 33 1 B2
rlabel metal1 84 35 84 35 1 Y
rlabel polysilicon 76 30 76 30 1 C1
rlabel polysilicon 36 57 36 57 1 A1
rlabel polysilicon 19 57 19 57 1 A2
rlabel polysilicon 53 57 53 57 1 B1
rlabel polysilicon 70 57 70 57 1 B1
<< end >>
