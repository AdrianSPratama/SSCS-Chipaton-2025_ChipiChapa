* SPICE3 file created from gf180mcu_gp9t3v3_oai221_1.2.ext - technology: gf180mcuD

.subckt gf180mcu_gp9t3v3_oai221_1 A0 A1 B0 B1 C Y vdd vss
X0 a_n110_n70# A1.t0 Y.t1 vss.t5 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X1 Y.t4 B1.t0 a_560_410# vdd.t7 pfet_03v3 ad=0.85p pd=4.4u as=0.2125p ps=1.95u w=1.7u l=0.3u
X2 a_390_n70# C.t0 a_n110_n70# vss.t6 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X3 a_390_n70# B1.t1 vss.t4 vss.t3 nfet_03v3 ad=0.425p pd=2.7u as=0.23375p ps=1.4u w=0.85u l=0.3u
X4 a_110_410# A0.t0 vdd.t1 vdd.t0 pfet_03v3 ad=0.2125p pd=1.95u as=0.85p ps=4.4u w=1.7u l=0.3u
X5 Y.t2 A1.t1 a_110_410# vdd.t4 pfet_03v3 ad=0.4675p pd=2.25u as=0.2125p ps=1.95u w=1.7u l=0.3u
X6 vss.t1 B0.t0 a_390_n70# vss.t0 nfet_03v3 ad=0.23375p pd=1.4u as=0.23375p ps=1.4u w=0.85u l=0.3u
X7 vdd.t6 C.t1 Y.t3 vdd.t5 pfet_03v3 ad=0.4675p pd=2.25u as=0.4675p ps=2.25u w=1.7u l=0.3u
X8 Y.t0 A0.t1 a_n110_n70# vss.t2 nfet_03v3 ad=0.23375p pd=1.4u as=0.425p ps=2.7u w=0.85u l=0.3u
X9 a_560_410# B0.t1 vdd.t3 vdd.t2 pfet_03v3 ad=0.2125p pd=1.95u as=0.4675p ps=2.25u w=1.7u l=0.3u
C0 vdd Y 0.50179f
C1 B1 a_390_n70# 0.1264f
C2 B1 B0 0.16085f
C3 B0 a_390_n70# 0.12515f
C4 vdd A0 0.15311f
C5 a_n110_n70# Y 0.15769f
C6 A1 Y 0.17058f
C7 C Y 0.14177f
C8 a_n110_n70# A0 0.05779f
C9 B1 vdd 0.12123f
C10 A1 A0 0.08267f
C11 vdd a_110_410# 0.00549f
C12 vdd a_390_n70# 0
C13 C A0 0
C14 vdd B0 0.0949f
C15 a_560_410# Y 0.00573f
C16 a_n110_n70# a_390_n70# 0.06353f
C17 a_n110_n70# B0 0
C18 B1 A1 0
C19 A1 a_390_n70# 0
C20 A1 B0 0.00127f
C21 C a_390_n70# 0.02952f
C22 C B0 0.1392f
C23 A0 Y 0.09132f
C24 B0 a_560_410# 0.00204f
C25 a_n110_n70# vdd 0.00585f
C26 A1 vdd 0.0909f
C27 C vdd 0.10899f
C28 B1 Y 0.14349f
C29 a_110_410# Y 0.00573f
C30 Y a_390_n70# 0.05423f
C31 B0 Y 0.13041f
C32 a_n110_n70# A1 0.05638f
C33 a_n110_n70# C 0.00479f
C34 vdd a_560_410# 0.00549f
C35 A1 C 0.10829f
R0 A1.n0 A1.t1 43.8005
R1 A1.n0 A1.t0 20.0755
R2 A1 A1.n0 12.5342
R3 Y.n2 Y.n1 7.0925
R4 Y.n5 Y.n4 4.5455
R5 Y.n3 Y.t4 3.24419
R6 Y.n2 Y.n0 2.12983
R7 Y.n1 Y.t1 2.03874
R8 Y.n1 Y.t0 2.03874
R9 Y.n0 Y.t3 1.13285
R10 Y.n0 Y.t2 1.13285
R11 Y.n3 Y.n2 0.8285
R12 Y Y.n5 0.03425
R13 Y.n5 Y 0.03425
R14 Y.n4 Y.n3 0.0305
R15 vss.t0 vss.t6 891.13
R16 vss.t5 vss.n7 864.919
R17 vss.n4 vss.t3 707.662
R18 vss.t2 vss.n8 655.242
R19 vss.n9 vss.t2 450.764
R20 vss.t3 vss.n3 403.649
R21 vss.n8 vss.t5 235.887
R22 vss.n4 vss.t0 183.469
R23 vss.n7 vss.t6 26.2102
R24 vss.n5 vss.n4 10.4005
R25 vss.n7 vss.n6 10.4005
R26 vss.n8 vss.n0 10.4005
R27 vss.n3 vss.n2 6.5885
R28 vss vss.n9 5.2005
R29 vss.n2 vss.t4 2.03874
R30 vss.n2 vss.t1 2.03874
R31 vss.n9 vss.n1 1.94494
R32 vss.n6 vss.n5 0.1355
R33 vss.n6 vss.n0 0.1355
R34 vss vss.n0 0.1355
R35 vss.n5 vss.n3 0.0326429
R36 B1.n0 B1.t0 40.1505
R37 B1.n0 B1.t1 23.7255
R38 B1 B1.n0 12.5342
R39 vdd.t5 vdd.t2 265.625
R40 vdd.n5 vdd.t4 257.812
R41 vdd.n9 vdd.t0 232.863
R42 vdd.t0 vdd.n8 101.562
R43 vdd.n4 vdd.t7 74.1583
R44 vdd.n8 vdd.t4 70.313
R45 vdd.t2 vdd.n4 58.866
R46 vdd.n6 vdd.n5 12.6005
R47 vdd.n8 vdd.n7 12.6005
R48 vdd.n4 vdd.n3 8.05153
R49 vdd.n5 vdd.t5 7.813
R50 vdd vdd.n9 6.3005
R51 vdd.n0 vdd.t1 3.29819
R52 vdd.n3 vdd.n2 2.16583
R53 vdd.n9 vdd.n1 1.7505
R54 vdd.n2 vdd.t3 1.13285
R55 vdd.n2 vdd.t6 1.13285
R56 vdd.n7 vdd.n6 0.1355
R57 vdd.n7 vdd.n0 0.0969286
R58 vdd.n6 vdd.n3 0.0583571
R59 vdd vdd.n0 0.0390714
R60 C.n0 C.t1 40.1505
R61 C.n0 C.t0 23.7255
R62 C C.n0 12.5342
R63 A0.n0 A0.t0 43.8005
R64 A0.n0 A0.t1 20.0755
R65 A0 A0.n0 12.5342
R66 B0.n0 B0.t1 40.1505
R67 B0.n0 B0.t0 23.7255
R68 B0 B0.n0 12.5342
C36 Y vss 0.28022f
C37 B1 vss 0.33834f
C38 B0 vss 0.25665f
C39 C vss 0.27627f
C40 A1 vss 0.28049f
C41 A0 vss 0.36107f
C42 vdd vss 2.36999f
C43 a_390_n70# vss 0.32897f 
C44 a_n110_n70# vss 0.49548f 
.ends